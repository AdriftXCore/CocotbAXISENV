`ifndef __TOP_DEFINE_VH
`define __TOP_DEFINE_VH 1

`define DATA_W 128

`endif